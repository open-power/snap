/afs/vlsilab.boeblingen.ibm.com/proj/fpga/framework/castella/snap_9V3_init/snap/hardware/hdl/core/dma_rams_capi20.vhd_source